
`include "sys_def.svh"
`include "ISA.svh"

module testbench;



endmodule
