`include "sys_defs.svh"

module load_queue (
    input logic clock, reset,
    
);

endmodule