`include "sys_defs.svh"

module prf #(
    parameter SIZE = `PHYS_REG_SZ_R10K
)(
    input clock, reset,
    
);

endmodule
