`include "sys_defs.svh"

module testbench;
    parameter SIZE = `ARCH_REG_SZ;

    logic clock, reset, correct;

    // input 
    RRAT_CT_INPUT rrat_ct_input;

    // output
    




endmodule;