`include "sys_defs.svh"
    
endtask

module ras #(
    parameter PORTS = `N,
    parameter DEPTH = 4
) (
    input clock, reset,

);
    
endmodule
